module counter_8bit (
    input  wire       clk,
    input  wire       reset,
    input  wire       enable,
    output reg  [7:0] count
);


endmodule
