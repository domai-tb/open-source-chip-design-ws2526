module barrel_shifter (
    input  wire [3:0] data_in,
    input  wire [2:0] shift_amt,
    input  wire       direction,
    output reg  [3:0] data_out
);


endmodule
