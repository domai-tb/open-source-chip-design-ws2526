module half_adder (
    input  wire a,
    input  wire b,
    output wire sum,
    output wire carry
);


endmodule